library ieee;
use ieee.std_logic_1164.all;

entity Keccak_parallel is
  port(
  clk:in std_logic);
end Keccak_parallel;

architecture beh of Keccak_parallel is
begin
end beh;